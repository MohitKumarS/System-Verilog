interface pif (input clk, rst);
  
endinterface
