class adder_tx;
  int a = 1;
  int b = 2;
  
  function print();
    $display("Printing Transaction :\n a = %0d \n b = %0d",a,b);
  endfunction
endclass
