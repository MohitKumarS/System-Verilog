class adder_gen;
  task run();
    $display("I'm in adder_gen");
  endtask
endclass
