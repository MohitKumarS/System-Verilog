class common;
  static mailbox gen2bfm = new();
  //static virtual intf vif;
endclass

