interface adder_intf (input clk, rst);
  logic [31:0] data;
  logic [31:0] addr;
  
endinterface
