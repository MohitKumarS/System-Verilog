class adder_bfm;
  task run();
    $display("I'm in adder_bfm");
  endtask
endclass
