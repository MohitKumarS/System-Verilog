
`include "adder_intf.sv"

`include "common.sv"

`include "adder_tx.sv"

`include "adder_gen.sv"

`include "adder_bfm.sv"

`include "adder_agent.sv"

`include "adder_env.sv"

`include "adder_test.sv"

`include "top.sv"

